module square_root_unit(
			reset,
			clk,
			e,
			f
			);

input 
      reset,
      clk;

input [30:0] e;   //31-bit input from log_unit block

output [16:0] f;  //17-bit output

//parameter C2_f = 0.54506876 ;
//parameter C1_f = 0.50332717 ;
//parameter C0_f = -0.03541023 ;

//parameter C2_f = 9144736;
//parameter C1_f = 8444428;
//parameter C0_f = -594085;

parameter C2_f = 40'h00008b899f;
parameter C1_f = 40'h000080da0c;
parameter C0_f = 40'hfffff6ef5a;

parameter SQ_SEL_BITS = 6;

wire [47:0] din;
wire [5:0] numz;

reg [6:0] exp_f;
reg [16:0] x_f_p;
reg [16:0] x_f;
reg signed [16:0] y_f_reg_1;
reg signed [16:0] y_f_reg_2;
reg [6:0] exp_f_p;
reg [16:0] f;

reg [11:0] coef1 ;
reg [19:0] coef0 ;

reg [11:0] coef1_reg ;
reg [19:0] coef0_reg ;

assign din = {e, 17'h1ffff};

lzd lzd (
              .reset(reset),
              .clk(clk),
              .din(din),
              .numz(numz)
	);

always @(posedge clk or posedge reset)
begin
if (reset)
        begin
        exp_f <= 0;
        x_f_p <= 0;
        exp_f_p <= 0;
        x_f <= 0;
        coef1_reg <= 0;
        coef0_reg <= 0;
        y_f_reg_1 <= 0;
        y_f_reg_2 <= 0;
        f <= 0;
        end
else
        begin
        // Range Reduction
        exp_f <= 5 - numz;
        x_f_p <= e >> exp_f;
        exp_f_p <= exp_f[0] ? (exp_f + 1) >> 1 : exp_f >> 1 ;
        x_f <= exp_f[0] ? x_f_p >> 1 : x_f_p ;
        coef1_reg <= coef1;
        coef0_reg <= coef0;

        y_f_reg_1 <= $signed(coef1_reg) * $signed(x_f[16-SQ_SEL_BITS:0]) ;
        y_f_reg_2 <= $signed(coef0_reg) * $signed(y_f_reg_1) ;

        // Range Reconstruction
        f <= y_f_reg_2 << exp_f_p ;
        end
end

// Square Root Coefficients

wire [SQ_SEL_BITS-1:0] sel = x_f[16:16-(SQ_SEL_BITS-1)] ;

always @(sel)
begin
  case(sel)
       0 : {coef1[11:0], coef0[19:0]} =   32'b000_011111101___000_10000001011101111;
       1 : {coef1[11:0], coef0[19:0]} =   32'b000_011110111___000_10000100011001101;
       2 : {coef1[11:0], coef0[19:0]} =   32'b000_011110010___000_10000111010001010;
       3 : {coef1[11:0], coef0[19:0]} =   32'b000_011101101___000_10001010000101001;
       4 : {coef1[11:0], coef0[19:0]} =   32'b000_011101001___000_10001100110101011;
       5 : {coef1[11:0], coef0[19:0]} =   32'b000_011100100___000_10001111100010011;
       6 : {coef1[11:0], coef0[19:0]} =   32'b000_011100000___000_10010010001100000;
       7 : {coef1[11:0], coef0[19:0]} =   32'b000_011011100___000_10010100110010101;
       8 : {coef1[11:0], coef0[19:0]} =   32'b000_011011000___000_10010111010110100;
       9 : {coef1[11:0], coef0[19:0]} =   32'b000_011010101___000_10011001110111100;
      10 : {coef1[11:0], coef0[19:0]} =   32'b000_011010010___000_10011100010110000;
      11 : {coef1[11:0], coef0[19:0]} =   32'b000_011001110___000_10011110110010000;
      12 : {coef1[11:0], coef0[19:0]} =   32'b000_011001011___000_10100001001011101;
      13 : {coef1[11:0], coef0[19:0]} =   32'b000_011001000___000_10100011100011000;
      14 : {coef1[11:0], coef0[19:0]} =   32'b000_011000110___000_10100101111000010;
      15 : {coef1[11:0], coef0[19:0]} =   32'b000_011000011___000_10101000001011100;
      16 : {coef1[11:0], coef0[19:0]} =   32'b000_011000000___000_10101010011100101;
      17 : {coef1[11:0], coef0[19:0]} =   32'b000_010111110___000_10101100101011111;
      18 : {coef1[11:0], coef0[19:0]} =   32'b000_010111011___000_10101110111001010;
      19 : {coef1[11:0], coef0[19:0]} =   32'b000_010111001___000_10110001000101000;
      20 : {coef1[11:0], coef0[19:0]} =   32'b000_010110111___000_10110011001110111;
      21 : {coef1[11:0], coef0[19:0]} =   32'b000_010110101___000_10110101010111010;
      22 : {coef1[11:0], coef0[19:0]} =   32'b000_010110011___000_10110111011110000;
      23 : {coef1[11:0], coef0[19:0]} =   32'b000_010110001___000_10111001100011010;
      24 : {coef1[11:0], coef0[19:0]} =   32'b000_010101111___000_10111011100110111;
      25 : {coef1[11:0], coef0[19:0]} =   32'b000_010101101___000_10111101101001010;
      26 : {coef1[11:0], coef0[19:0]} =   32'b000_010101011___000_10111111101010001;
      27 : {coef1[11:0], coef0[19:0]} =   32'b000_010101001___000_11000001101001110;
      28 : {coef1[11:0], coef0[19:0]} =   32'b000_010101000___000_11000011101000000;
      29 : {coef1[11:0], coef0[19:0]} =   32'b000_010100110___000_11000101100101000;
      30 : {coef1[11:0], coef0[19:0]} =   32'b000_010100100___000_11000111100000110;
      31 : {coef1[11:0], coef0[19:0]} =   32'b000_010100011___000_11001001011011011;
      32 : {coef1[11:0], coef0[19:0]} =   32'b000_010100001___000_11001011010100111;
      33 : {coef1[11:0], coef0[19:0]} =   32'b000_010100000___000_11001101001101001;
      34 : {coef1[11:0], coef0[19:0]} =   32'b000_010011110___000_11001111000100011;
      35 : {coef1[11:0], coef0[19:0]} =   32'b000_010011101___000_11010000111010100;
      36 : {coef1[11:0], coef0[19:0]} =   32'b000_010011011___000_11010010101111110;
      37 : {coef1[11:0], coef0[19:0]} =   32'b000_010011010___000_11010100100011110;
      38 : {coef1[11:0], coef0[19:0]} =   32'b000_010011001___000_11010110010111000;
      39 : {coef1[11:0], coef0[19:0]} =   32'b000_010011000___000_11011000001001001;
      40 : {coef1[11:0], coef0[19:0]} =   32'b000_010010110___000_11011001111010011;
      41 : {coef1[11:0], coef0[19:0]} =   32'b000_010010101___000_11011011101010110;
      42 : {coef1[11:0], coef0[19:0]} =   32'b000_010010100___000_11011101011010001;
      43 : {coef1[11:0], coef0[19:0]} =   32'b000_010010011___000_11011111001000110;
      44 : {coef1[11:0], coef0[19:0]} =   32'b000_010010010___000_11100000110110100;
      45 : {coef1[11:0], coef0[19:0]} =   32'b000_010010001___000_11100010100011011;
      46 : {coef1[11:0], coef0[19:0]} =   32'b000_010010000___000_11100100001111011;
      47 : {coef1[11:0], coef0[19:0]} =   32'b000_010001111___000_11100101111010110;
      48 : {coef1[11:0], coef0[19:0]} =   32'b000_010001101___000_11100111100101010;
      49 : {coef1[11:0], coef0[19:0]} =   32'b000_010001100___000_11101001001111000;
      50 : {coef1[11:0], coef0[19:0]} =   32'b000_010001100___000_11101010111000000;
      51 : {coef1[11:0], coef0[19:0]} =   32'b000_010001011___000_11101100100000010;
      52 : {coef1[11:0], coef0[19:0]} =   32'b000_010001010___000_11101110000111110;
      53 : {coef1[11:0], coef0[19:0]} =   32'b000_010001001___000_11101111101110101;
      54 : {coef1[11:0], coef0[19:0]} =   32'b000_010001000___000_11110001010100111;
      55 : {coef1[11:0], coef0[19:0]} =   32'b000_010000111___000_11110010111010011;
      56 : {coef1[11:0], coef0[19:0]} =   32'b000_010000110___000_11110100011111010;
      57 : {coef1[11:0], coef0[19:0]} =   32'b000_010000101___000_11110110000011011;
      58 : {coef1[11:0], coef0[19:0]} =   32'b000_010000100___000_11110111100111000;
      59 : {coef1[11:0], coef0[19:0]} =   32'b000_010000100___000_11111001001001111;
      60 : {coef1[11:0], coef0[19:0]} =   32'b000_010000011___000_11111010101100010;
      61 : {coef1[11:0], coef0[19:0]} =   32'b000_010000010___000_11111100001110000;
      62 : {coef1[11:0], coef0[19:0]} =   32'b000_010000001___000_11111101101111001;
      63 : {coef1[11:0], coef0[19:0]} =   32'b000_010000000___000_11111111001111110;
  endcase
end

endmodule
