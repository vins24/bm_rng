module log_unit (
		 reset,
	         clk,
		 u0,
		 e
		);

input reset,
      clk;

input [47:0] u0;

output [30:0] e;     //e(31,24) 

//parameter C2_e = 1.14458115 ;
//parameter C1_e = -1.38438915 ;
//parameter C0_e = 0.23388019 ;
//parameter ln2 = 0.69314718;

//parameter C2_e = 19202884;
//parameter C1_e = -23226194;
//parameter C0_e = 3923858;
//parameter ln2 = 11629079;

parameter C2_e = 40'h0001250344;
parameter C1_e = 40'hfffe9d98ad;
parameter C0_e = 40'h00003bdf92;
parameter ln2 =  40'h0000b17217;
parameter LN_SEL_BITS =  8;

wire [47:0] u0;
wire [5:0] numz;

reg [6:0] exp_e;
reg [47:0] x_e;
reg signed [30:0] e_p;

reg signed [30:0] y_e_reg_1;
reg signed [30:0] y_e_reg_2;
reg signed [30:0] y_e_reg_3;
reg signed [30:0] y_e_reg_4;

reg signed [12:0] coef2 ;
reg signed [21:0] coef1 ;
reg signed [29:0] coef0 ;
reg signed [30:0] e_pp;
reg signed [30:0] e;

lzd lzd (
              .reset(reset),
              .clk(clk),
              .din(u0),
              .numz(numz)
             );

always @(posedge clk or posedge reset)
begin
if (reset)
        begin
        exp_e <= 0;
        x_e <= 0;
	e_p <= 0;
        y_e_reg_1 <= 0;
        y_e_reg_2 <= 0;
        y_e_reg_3 <= 0;
        y_e_reg_4 <= 0;
        y_e_reg_4 <= 0;
        e_pp <= 0;
        e <= 0;
        end
else
        begin
        // Range Reduction
        exp_e <= numz + 1;
        x_e <= u0 << exp_e;

	e_p <= $signed(exp_e) * $signed(ln2);

        y_e_reg_1 <= $signed(coef2) * $signed(x_e[30-LN_SEL_BITS:0]) ;
        y_e_reg_2 <= $signed(coef1) + $signed(y_e_reg_1) ;
        y_e_reg_3 <= $signed(x_e[30-LN_SEL_BITS:0]) * $signed(y_e_reg_2) ;
        y_e_reg_4 <= $signed(coef0) + $signed(y_e_reg_3) ;
        // Range Reconstruction
        e_pp <= $signed(e_p) - $signed(y_e_reg_1);
        e <= e_pp << 1;
        end
end

// Natural Log Coefficients

wire [LN_SEL_BITS-1:0] sel = x_e[30:30-(LN_SEL_BITS-1)] ;

always @(sel)
begin
  case(sel)
       0 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0000001000___000_1111111100000101010___111_111111110000000110000000000;
       1 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0000010000___000_1111111000001001001___111_111111100000001111111000000;
       2 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0000010111___000_1111110100001111000___111_111111010000011101110000000;
       3 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0000011111___000_1111110000010110110___111_111111000000101111100000000;
       4 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0000100111___000_1111101100100000011___111_111110110001000101000000000;
       5 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0000101110___000_1111101000101011111___111_111110100001011110011000000;
       6 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0000110110___000_1111100100111001010___111_111110010001111011100000000;
       7 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0000111101___000_1111100001001000100___111_111110000010011100100000000;
       8 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0001000100___000_1111011101011001100___111_111101110011000001001000000;
       9 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0001001011___000_1111011001101100011___111_111101100011101001100000000;
      10 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0001010010___000_1111010110000000111___111_111101010100010101100000000;
      11 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0001011001___000_1111010010010111010___111_111101000101000101010000000;
      12 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0001100000___000_1111001110101111010___111_111100110101111000100000000;
      13 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0001100111___000_1111001011001001001___111_111100100110101111011000000;
      14 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0001101110___000_1111000111100100100___111_111100010111101001111000000;
      15 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0001110100___000_1111000100000001110___111_111100001000100111111000000;
      16 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0001111011___000_1111000000100000100___111_111011111001101001100000000;
      17 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0010000010___000_1110111101000000111___111_111011101010101110100000000;
      18 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0010001000___000_1110111001100011000___111_111011011011110111000000000;
      19 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0010001111___000_1110110110000110101___111_111011001101000010111000000;
      20 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0010010101___000_1110110010101011111___111_111010111110010010010000000;
      21 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0010011011___000_1110101111010010110___111_111010101111100101000000000;
      22 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0010100001___000_1110101011111011001___111_111010100000111011001000000;
      23 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0010100111___000_1110101000100101000___111_111010010010010100100000000;
      24 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0010101101___000_1110100101010000011___111_111010000011110001010000000;
      25 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0010110011___000_1110100001111101011___111_111001110101010001011000000;
      26 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0010111001___000_1110011110101011110___111_111001100110110100110000000;
      27 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0010111111___000_1110011011011011101___111_111001011000011011010000000;
      28 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0011000101___000_1110011000001101000___111_111001001010000101001000000;
      29 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0011001011___000_1110010100111111110___111_111000111011110010001000000;
      30 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0011010001___000_1110010001110011111___111_111000101101100010011000000;
      31 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0011010110___000_1110001110101001100___111_111000011111010101110000000;
      32 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0011011100___000_1110001011100000100___111_111000010001001100010000000;
      33 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0011100001___000_1110001000011001000___111_111000000011000101110000000;
      34 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0011100111___000_1110000101010010110___111_110111110101000010100000000;
      35 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0011101100___000_1110000010001101111___111_110111100111000010010000000;
      36 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0011110010___000_1101111111001010010___111_110111011001000101001000000;
      37 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0011110111___000_1101111100001000000___111_110111001011001011000000000;
      38 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0011111100___000_1101111001000111001___111_110110111101010011111000000;
      39 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0100000001___000_1101110110000111100___111_110110101111011111110000000;
      40 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0100000110___000_1101110011001001010___111_110110100001101110101000000;
      41 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0100001011___000_1101110000001100001___111_110110010100000000011000000;
      42 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0100010000___000_1101101101010000011___111_110110000110010101001000000;
      43 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0100010101___000_1101101010010101111___111_110101111000101100110000000;
      44 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0100011010___000_1101100111011100100___111_110101101011000111011000000;
      45 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0100011111___000_1101100100100100100___111_110101011101100100110000000;
      46 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0100100100___000_1101100001101101101___111_110101010000000101000000000;
      47 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0100101001___000_1101011110110111111___111_110101000010101000001000000;
      48 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0100101110___000_1101011100000011011___111_110100110101001110000000000;
      49 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0100110010___000_1101011001010000001___111_110100100111110110110000000;
      50 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0100110111___000_1101010110011110000___111_110100011010100010010000000;
      51 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0100111100___000_1101010011101101000___111_110100001101010000100000000;
      52 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101000000___000_1101010000111101001___111_110100000000000001100000000;
      53 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101000101___000_1101001110001110011___111_110011110010110101010000000;
      54 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101001001___000_1101001011100000110___111_110011100101101011110000000;
      55 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101001110___000_1101001000110100011___111_110011011000100100111000000;
      56 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101010010___000_1101000110001000111___111_110011001011100000110000000;
      57 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101010110___000_1101000011011110101___111_110010111110011111001000000;
      58 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101011011___000_1101000000110101011___111_110010110001100000010000000;
      59 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101011111___000_1100111110001101010___111_110010100100100100000000000;
      60 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101100011___000_1100111011100110001___111_110010010111101010011000000;
      61 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101100111___000_1100111001000000001___111_110010001010110011011000000;
      62 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101101011___000_1100110110011011001___111_110001111101111110111000000;
      63 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101110000___000_1100110011110111001___111_110001110001001100111000000;
      64 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101110100___000_1100110001010100001___111_110001100100011101100000000;
      65 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101111000___000_1100101110110010001___111_110001010111110000110000000;
      66 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0101111100___000_1100101100010001010___111_110001001011000110011000000;
      67 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110000000___000_1100101001110001010___111_110000111110011110100000000;
      68 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110000100___000_1100100111010010010___111_110000110001111001001000000;
      69 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110000111___000_1100100100110100010___111_110000100101010110010000000;
      70 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110001011___000_1100100010010111010___111_110000011000110101111000000;
      71 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110001111___000_1100011111111011001___111_110000001100010111111000000;
      72 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110010011___000_1100011101100000000___111_101111111111111100010000000;
      73 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110010111___000_1100011011000101110___111_101111110011100011001000000;
      74 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110011010___000_1100011000101100100___111_101111100111001100010000000;
      75 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110011110___000_1100010110010100001___111_101111011010110111111000000;
      76 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110100010___000_1100010011111100101___111_101111001110100101111000000;
      77 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110100101___000_1100010001100110001___111_101111000010010110001000000;
      78 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110101001___000_1100001111010000100___111_101110110110001000110000000;
      79 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110101100___000_1100001100111011110___111_101110101001111101110000000;
      80 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110110000___000_1100001010100111111___111_101110011101110101000000000;
      81 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110110011___000_1100001000010100111___111_101110010001101110101000000;
      82 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110110111___000_1100000110000010110___111_101110000101101010100000000;
      83 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110111010___000_1100000011110001011___111_101101111001101000101000000;
      84 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0110111110___000_1100000001100001000___111_101101101101101001000000000;
      85 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111000001___000_1011111111010001011___111_101101100001101011101000000;
      86 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111000100___000_1011111101000010101___111_101101010101110000011000000;
      87 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111001000___000_1011111010110100110___111_101101001001110111100000000;
      88 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111001011___000_1011111000100111101___111_101100111110000000110000000;
      89 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111001110___000_1011110110011011011___111_101100110010001100010000000;
      90 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111010010___000_1011110100001111111___111_101100100110011001111000000;
      91 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111010101___000_1011110010000101001___111_101100011010101001101000000;
      92 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111011000___000_1011101111111011010___111_101100001110111011100000000;
      93 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111011011___000_1011101101110010001___111_101100000011001111101000000;
      94 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111011110___000_1011101011101001110___111_101011110111100101111000000;
      95 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111100001___000_1011101001100010010___111_101011101011111110010000000;
      96 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111100100___000_1011100111011011100___111_101011100000011000101000000;
      97 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111100111___000_1011100101010101011___111_101011010100110101001000000;
      98 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111101010___000_1011100011010000001___111_101011001001010011110000000;
      99 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111101101___000_1011100001001011101___111_101010111101110100011000000;
     100 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111110000___000_1011011111000111110___111_101010110010010111001000000;
     101 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111110011___000_1011011101000100110___111_101010100110111011111000000;
     102 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111110110___000_1011011011000010011___111_101010011011100010110000000;
     103 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111111001___000_1011011001000000110___111_101010010000001011100000000;
     104 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111111100___000_1011010110111111111___111_101010000100110110011000000;
     105 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_0111111111___000_1011010100111111110___111_101001111001100011010000000;
     106 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000000010___000_1011010011000000010___111_101001101110010010001000000;
     107 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000000100___000_1011010001000001100___111_101001100011000010111000000;
     108 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000000111___000_1011001111000011011___111_101001010111110101101000000;
     109 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000001010___000_1011001101000110000___111_101001001100101010011000000;
     110 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000001101___000_1011001011001001010___111_101001000001100001001000000;
     111 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000001111___000_1011001001001101010___111_101000110110011001110000000;
     112 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000010010___000_1011000111010001111___111_101000101011010100010000000;
     113 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000010101___000_1011000101010111001___111_101000100000010000110000000;
     114 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000010111___000_1011000011011101001___111_101000010101001111001000000;
     115 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000011010___000_1011000001100011110___111_101000001010001111011000000;
     116 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000011100___000_1010111111101011000___111_100111111111010001100000000;
     117 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000011111___000_1010111101110010111___111_100111110100010101100000000;
     118 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000100010___000_1010111011111011011___111_100111101001011011011000000;
     119 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000100100___000_1010111010000100101___111_100111011110100011001000000;
     120 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000100111___000_1010111000001110011___111_100111010011101100101000000;
     121 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000101001___000_1010110110011000111___111_100111001000111000001000000;
     122 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000101100___000_1010110100100011111___111_100110111110000101011000000;
     123 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000101110___000_1010110010101111100___111_100110110011010100011000000;
     124 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000110001___000_1010110000111011110___111_100110101000100101010000000;
     125 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000110011___000_1010101111001000101___111_100110011101110111111000000;
     126 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000110101___000_1010101101010110001___111_100110010011001100011000000;
     127 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000111000___000_1010101011100100010___111_100110001000100010100000000;
     128 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000111010___000_1010101001110010111___111_100101111101111010100000000;
     129 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000111100___000_1010101000000010001___111_100101110011010100010000000;
     130 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1000111111___000_1010100110010001111___111_100101101000101111110000000;
     131 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001000001___000_1010100100100010011___111_100101011110001101000000000;
     132 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001000011___000_1010100010110011010___111_100101010011101100000000000;
     133 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001000110___000_1010100001000100111___111_100101001001001100101000000;
     134 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001001000___000_1010011111010111000___111_100100111110101111001000000;
     135 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001001010___000_1010011101101001101___111_100100110100010011010000000;
     136 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001001100___000_1010011011111100111___111_100100101001111001000000000;
     137 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001001111___000_1010011010010000101___111_100100011111100000100000000;
     138 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001010001___000_1010011000100100111___111_100100010101001001110000000;
     139 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001010011___000_1010010110111001110___111_100100001010110100100000000;
     140 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001010101___000_1010010101001111010___111_100100000000100001001000000;
     141 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001010111___000_1010010011100101001___111_100011110110001111010000000;
     142 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001011001___000_1010010001111011101___111_100011101011111111000000000;
     143 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001011011___000_1010010000010010101___111_100011100001110000100000000;
     144 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001011101___000_1010001110101010001___111_100011010111100011101000000;
     145 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001100000___000_1010001101000010001___111_100011001101011000010000000;
     146 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001100010___000_1010001011011010101___111_100011000011001110101000000;
     147 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001100100___000_1010001001110011110___111_100010111001000110101000000;
     148 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001100110___000_1010001000001101010___111_100010101111000000001000000;
     149 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001101000___000_1010000110100111011___111_100010100100111011010000000;
     150 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001101010___000_1010000101000001111___111_100010011010110111111000000;
     151 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001101100___000_1010000011011101000___111_100010010000110110010000000;
     152 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001101110___000_1010000001111000100___111_100010000110110110000000000;
     153 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001110000___000_1010000000010100101___111_100001111100110111011000000;
     154 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001110010___000_1001111110110001001___111_100001110010111010011000000;
     155 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001110011___000_1001111101001110001___111_100001101000111110111000000;
     156 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001110101___000_1001111011101011101___111_100001011111000100111000000;
     157 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001110111___000_1001111010001001101___111_100001010101001100100000000;
     158 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001111001___000_1001111000101000000___111_100001001011010101100000000;
     159 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001111011___000_1001110111000110111___111_100001000001100000001000000;
     160 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001111101___000_1001110101100110010___111_100000110111101100010000000;
     161 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1001111111___000_1001110100000110001___111_100000101101111001111000000;
     162 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010000001___000_1001110010100110011___111_100000100100001001000000000;
     163 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010000010___000_1001110001000111001___111_100000011010011001101000000;
     164 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010000100___000_1001101111101000011___111_100000010000101011101000000;
     165 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010000110___000_1001101110001010000___111_100000000110111111001000000;
     166 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010001000___000_1001101100101100000___111_011111111101010100010000000;
     167 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010001010___000_1001101011001110101___111_011111110011101010101000000;
     168 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010001011___000_1001101001110001100___111_011111101010000010100000000;
     169 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010001101___000_1001101000010101000___111_011111100000011011111000000;
     170 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010001111___000_1001100110111000110___111_011111010110110110110000000;
     171 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010010001___000_1001100101011101000___111_011111001101010011000000000;
     172 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010010010___000_1001100100000001110___111_011111000011110000101000000;
     173 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010010100___000_1001100010100110111___111_011110111010001111101000000;
     174 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010010110___000_1001100001001100011___111_011110110000110000001000000;
     175 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010010111___000_1001011111110010011___111_011110100111010010000000000;
     176 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010011001___000_1001011110011000110___111_011110011101110101010000000;
     177 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010011011___000_1001011100111111100___111_011110010100011010000000000;
     178 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010011100___000_1001011011100110110___111_011110001011000000000000000;
     179 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010011110___000_1001011010001110010___111_011110000001100111100000000;
     180 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010011111___000_1001011000110110010___111_011101111000010000010000000;
     181 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010100001___000_1001010111011110110___111_011101101110111010100000000;
     182 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010100011___000_1001010110000111100___111_011101100101100110000000000;
     183 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010100100___000_1001010100110000110___111_011101011100010010111000000;
     184 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010100110___000_1001010011011010010___111_011101010011000001001000000;
     185 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010100111___000_1001010010000100010___111_011101001001110000110000000;
     186 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010101001___000_1001010000101110101___111_011101000000100001101000000;
     187 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010101010___000_1001001111011001011___111_011100110111010011111000000;
     188 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010101100___000_1001001110000100100___111_011100101110000111100000000;
     189 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010101110___000_1001001100110000000___111_011100100100111100011000000;
     190 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010101111___000_1001001011011011111___111_011100011011110010100000000;
     191 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010110001___000_1001001010001000001___111_011100010010101010000000000;
     192 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010110010___000_1001001000110100111___111_011100001001100010111000000;
     193 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010110011___000_1001000111100001111___111_011100000000011101000000000;
     194 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010110101___000_1001000110001111010___111_011011110111011000011000000;
     195 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010110110___000_1001000100111101000___111_011011101110010101000000000;
     196 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010111000___000_1001000011101011000___111_011011100101010011000000000;
     197 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010111001___000_1001000010011001100___111_011011011100010010010000000;
     198 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010111011___000_1001000001001000011___111_011011010011010010110000000;
     199 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010111100___000_1000111111110111100___111_011011001010010100100000000;
     200 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010111110___000_1000111110100111000___111_011011000001010111100000000;
     201 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1010111111___000_1000111101010110111___111_011010111000011011110000000;
     202 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011000000___000_1000111100000111001___111_011010101111100001010000000;
     203 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011000010___000_1000111010110111110___111_011010100110101000000000000;
     204 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011000011___000_1000111001101000101___111_011010011101110000000000000;
     205 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011000100___000_1000111000011001111___111_011010010100111001001000000;
     206 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011000110___000_1000110111001011100___111_011010001100000011100000000;
     207 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011000111___000_1000110101111101011___111_011010000011001111010000000;
     208 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011001001___000_1000110100101111101___111_011001111010011100000000000;
     209 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011001010___000_1000110011100010010___111_011001110001101010001000000;
     210 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011001011___000_1000110010010101010___111_011001101000111001011000000;
     211 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011001101___000_1000110001001000100___111_011001100000001001111000000;
     212 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011001110___000_1000101111111100001___111_011001010111011011100000000;
     213 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011001111___000_1000101110110000000___111_011001001110101110011000000;
     214 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011010000___000_1000101101100100010___111_011001000110000010011000000;
     215 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011010010___000_1000101100011000110___111_011000111101010111100000000;
     216 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011010011___000_1000101011001101101___111_011000110100101101111000000;
     217 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011010100___000_1000101010000010111___111_011000101100000101100000000;
     218 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011010101___000_1000101000111000011___111_011000100011011110001000000;
     219 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011010111___000_1000100111101110001___111_011000011010111000000000000;
     220 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011011000___000_1000100110100100010___111_011000010010010011000000000;
     221 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011011001___000_1000100101011010110___111_011000001001101111001000000;
     222 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011011010___000_1000100100010001100___111_011000000001001100100000000;
     223 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011011100___000_1000100011001000100___111_010111111000101010111000000;
     224 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011011101___000_1000100001111111111___111_010111110000001010100000000;
     225 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011011110___000_1000100000110111100___111_010111100111101011001000000;
     226 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011011111___000_1000011111101111100___111_010111011111001101000000000;
     227 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011100000___000_1000011110100111110___111_010111010110101111111000000;
     228 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011100010___000_1000011101100000010___111_010111001110010100000000000;
     229 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011100011___000_1000011100011001001___111_010111000101111001001000000;
     230 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011100100___000_1000011011010010010___111_010110111101011111011000000;
     231 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011100101___000_1000011010001011101___111_010110110101000110110000000;
     232 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011100110___000_1000011001000101011___111_010110101100101111010000000;
     233 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011100111___000_1000010111111111011___111_010110100100011000110000000;
     234 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011101001___000_1000010110111001101___111_010110011100000011011000000;
     235 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011101010___000_1000010101110100001___111_010110010011101111001000000;
     236 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011101011___000_1000010100101111000___111_010110001011011100000000000;
     237 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011101100___000_1000010011101010001___111_010110000011001001110000000;
     238 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011101101___000_1000010010100101100___111_010101111010111000110000000;
     239 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011101110___000_1000010001100001010___111_010101110010101000110000000;
     240 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011101111___000_1000010000011101001___111_010101101010011001111000000;
     241 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011110000___000_1000001111011001011___111_010101100010001100000000000;
     242 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011110001___000_1000001110010101111___111_010101011001111111001000000;
     243 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011110011___000_1000001101010010101___111_010101010001110011011000000;
     244 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011110100___000_1000001100001111101___111_010101001001101000110000000;
     245 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011110101___000_1000001011001101000___111_010101000001011111000000000;
     246 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011110110___000_1000001010001010100___111_010100111001010110011000000;
     247 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011110111___000_1000001001001000011___111_010100110001001110110000000;
     248 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011111000___000_1000001000000110011___111_010100101001001000001000000;
     249 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011111001___000_1000000111000100110___111_010100100001000010101000000;
     250 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011111010___000_1000000110000011011___111_010100011000111110000000000;
     251 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011111011___000_1000000101000010010___111_010100010000111010100000000;
     252 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011111100___000_1000000100000001011___111_010100001000111000000000000;
     253 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011111101___000_1000000011000000110___111_010100000000110110100000000;
     254 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011111110___000_1000000010000000011___111_010011111000110110000000000;
     255 : {coef2[12:0], coef1[21:0], coef0[29:0]} =   65'b111_1011111111___000_1000000001000000010___111_010011110000110110100000000;
  endcase
end

endmodule 
