
module sin_cos_coef (
		     sel,
		     coef1,
		     coef0
		     );

input [6:0] sel;

output [11:0] coef1; 
output [18:0] coef0; 

// Cosine Coefficients

reg [11:0] coef1 ;
reg [18:0] coef0 ;

always @(sel)
begin
  case(sel)
       0 : {coef1[11:0], coef0[18:0]} =   31'b111_111111011___001_0000000000000000;
       1 : {coef1[11:0], coef0[18:0]} =   31'b111_111110001___001_0000000000001010;
       2 : {coef1[11:0], coef0[18:0]} =   31'b111_111100111___001_0000000000011110;
       3 : {coef1[11:0], coef0[18:0]} =   31'b111_111011101___001_0000000000111011;
       4 : {coef1[11:0], coef0[18:0]} =   31'b111_111010100___001_0000000001100011;
       5 : {coef1[11:0], coef0[18:0]} =   31'b111_111001010___001_0000000010010100;
       6 : {coef1[11:0], coef0[18:0]} =   31'b111_111000000___001_0000000011001111;
       7 : {coef1[11:0], coef0[18:0]} =   31'b111_110110110___001_0000000100010100;
       8 : {coef1[11:0], coef0[18:0]} =   31'b111_110101100___001_0000000101100010;
       9 : {coef1[11:0], coef0[18:0]} =   31'b111_110100010___001_0000000110111011;
      10 : {coef1[11:0], coef0[18:0]} =   31'b111_110011001___001_0000001000011101;
      11 : {coef1[11:0], coef0[18:0]} =   31'b111_110001111___001_0000001010001000;
      12 : {coef1[11:0], coef0[18:0]} =   31'b111_110000101___001_0000001011111101;
      13 : {coef1[11:0], coef0[18:0]} =   31'b111_101111011___001_0000001101111100;
      14 : {coef1[11:0], coef0[18:0]} =   31'b111_101110010___001_0000010000000100;
      15 : {coef1[11:0], coef0[18:0]} =   31'b111_101101000___001_0000010010010110;
      16 : {coef1[11:0], coef0[18:0]} =   31'b111_101011110___001_0000010100110000;
      17 : {coef1[11:0], coef0[18:0]} =   31'b111_101010101___001_0000010111010101;
      18 : {coef1[11:0], coef0[18:0]} =   31'b111_101001011___001_0000011010000010;
      19 : {coef1[11:0], coef0[18:0]} =   31'b111_101000001___001_0000011100111000;
      20 : {coef1[11:0], coef0[18:0]} =   31'b111_100111000___001_0000011111111000;
      21 : {coef1[11:0], coef0[18:0]} =   31'b111_100101110___001_0000100011000000;
      22 : {coef1[11:0], coef0[18:0]} =   31'b111_100100101___001_0000100110010001;
      23 : {coef1[11:0], coef0[18:0]} =   31'b111_100011011___001_0000101001101011;
      24 : {coef1[11:0], coef0[18:0]} =   31'b111_100010010___001_0000101101001110;
      25 : {coef1[11:0], coef0[18:0]} =   31'b111_100001000___001_0000110000111001;
      26 : {coef1[11:0], coef0[18:0]} =   31'b111_011111111___001_0000110100101101;
      27 : {coef1[11:0], coef0[18:0]} =   31'b111_011110110___001_0000111000101001;
      28 : {coef1[11:0], coef0[18:0]} =   31'b111_011101100___001_0000111100101101;
      29 : {coef1[11:0], coef0[18:0]} =   31'b111_011100011___001_0001000000111001;
      30 : {coef1[11:0], coef0[18:0]} =   31'b111_011011010___001_0001000101001101;
      31 : {coef1[11:0], coef0[18:0]} =   31'b111_011010001___001_0001001001101001;
      32 : {coef1[11:0], coef0[18:0]} =   31'b111_011001000___001_0001001110001101;
      33 : {coef1[11:0], coef0[18:0]} =   31'b111_010111111___001_0001010010111000;
      34 : {coef1[11:0], coef0[18:0]} =   31'b111_010110110___001_0001010111101011;
      35 : {coef1[11:0], coef0[18:0]} =   31'b111_010101101___001_0001011100100101;
      36 : {coef1[11:0], coef0[18:0]} =   31'b111_010100100___001_0001100001100110;
      37 : {coef1[11:0], coef0[18:0]} =   31'b111_010011011___001_0001100110101111;
      38 : {coef1[11:0], coef0[18:0]} =   31'b111_010010010___001_0001101011111101;
      39 : {coef1[11:0], coef0[18:0]} =   31'b111_010001001___001_0001110001010011;
      40 : {coef1[11:0], coef0[18:0]} =   31'b111_010000001___001_0001110110101111;
      41 : {coef1[11:0], coef0[18:0]} =   31'b111_001111000___001_0001111100010010;
      42 : {coef1[11:0], coef0[18:0]} =   31'b111_001101111___001_0010000001111010;
      43 : {coef1[11:0], coef0[18:0]} =   31'b111_001100111___001_0010000111101001;
      44 : {coef1[11:0], coef0[18:0]} =   31'b111_001011110___001_0010001101011101;
      45 : {coef1[11:0], coef0[18:0]} =   31'b111_001010110___001_0010010011010111;
      46 : {coef1[11:0], coef0[18:0]} =   31'b111_001001110___001_0010011001010111;
      47 : {coef1[11:0], coef0[18:0]} =   31'b111_001000101___001_0010011111011100;
      48 : {coef1[11:0], coef0[18:0]} =   31'b111_000111101___001_0010100101100110;
      49 : {coef1[11:0], coef0[18:0]} =   31'b111_000110101___001_0010101011110100;
      50 : {coef1[11:0], coef0[18:0]} =   31'b111_000101101___001_0010110010001000;
      51 : {coef1[11:0], coef0[18:0]} =   31'b111_000100101___001_0010111000100000;
      52 : {coef1[11:0], coef0[18:0]} =   31'b111_000011101___001_0010111110111100;
      53 : {coef1[11:0], coef0[18:0]} =   31'b111_000010101___001_0011000101011100;
      54 : {coef1[11:0], coef0[18:0]} =   31'b111_000001101___001_0011001100000000;
      55 : {coef1[11:0], coef0[18:0]} =   31'b111_000000110___001_0011010010101000;
      56 : {coef1[11:0], coef0[18:0]} =   31'b110_111111110___001_0011011001010011;
      57 : {coef1[11:0], coef0[18:0]} =   31'b110_111110110___001_0011100000000010;
      58 : {coef1[11:0], coef0[18:0]} =   31'b110_111101111___001_0011100110110011;
      59 : {coef1[11:0], coef0[18:0]} =   31'b110_111101000___001_0011101101100111;
      60 : {coef1[11:0], coef0[18:0]} =   31'b110_111100000___001_0011110100011110;
      61 : {coef1[11:0], coef0[18:0]} =   31'b110_111011001___001_0011111011010111;
      62 : {coef1[11:0], coef0[18:0]} =   31'b110_111010010___001_0100000010010010;
      63 : {coef1[11:0], coef0[18:0]} =   31'b110_111001011___001_0100001001001111;
      64 : {coef1[11:0], coef0[18:0]} =   31'b110_111000100___001_0100010000001110;
      65 : {coef1[11:0], coef0[18:0]} =   31'b110_110111101___001_0100010111001110;
      66 : {coef1[11:0], coef0[18:0]} =   31'b110_110110110___001_0100011110001111;
      67 : {coef1[11:0], coef0[18:0]} =   31'b110_110101111___001_0100100101010001;
      68 : {coef1[11:0], coef0[18:0]} =   31'b110_110101001___001_0100101100010100;
      69 : {coef1[11:0], coef0[18:0]} =   31'b110_110100010___001_0100110011010111;
      70 : {coef1[11:0], coef0[18:0]} =   31'b110_110011100___001_0100111010011010;
      71 : {coef1[11:0], coef0[18:0]} =   31'b110_110010101___001_0101000001011101;
      72 : {coef1[11:0], coef0[18:0]} =   31'b110_110001111___001_0101001000100000;
      73 : {coef1[11:0], coef0[18:0]} =   31'b110_110001001___001_0101001111100010;
      74 : {coef1[11:0], coef0[18:0]} =   31'b110_110000011___001_0101010110100011;
      75 : {coef1[11:0], coef0[18:0]} =   31'b110_101111101___001_0101011101100011;
      76 : {coef1[11:0], coef0[18:0]} =   31'b110_101110111___001_0101100100100010;
      77 : {coef1[11:0], coef0[18:0]} =   31'b110_101110001___001_0101101011011111;
      78 : {coef1[11:0], coef0[18:0]} =   31'b110_101101100___001_0101110010011011;
      79 : {coef1[11:0], coef0[18:0]} =   31'b110_101100110___001_0101111001010100;
      80 : {coef1[11:0], coef0[18:0]} =   31'b110_101100001___001_0110000000001010;
      81 : {coef1[11:0], coef0[18:0]} =   31'b110_101011011___001_0110000110111110;
      82 : {coef1[11:0], coef0[18:0]} =   31'b110_101010110___001_0110001101101111;
      83 : {coef1[11:0], coef0[18:0]} =   31'b110_101010001___001_0110010100011101;
      84 : {coef1[11:0], coef0[18:0]} =   31'b110_101001100___001_0110011011000111;
      85 : {coef1[11:0], coef0[18:0]} =   31'b110_101000111___001_0110100001101110;
      86 : {coef1[11:0], coef0[18:0]} =   31'b110_101000010___001_0110101000010000;
      87 : {coef1[11:0], coef0[18:0]} =   31'b110_100111101___001_0110101110101110;
      88 : {coef1[11:0], coef0[18:0]} =   31'b110_100111000___001_0110110101000111;
      89 : {coef1[11:0], coef0[18:0]} =   31'b110_100110100___001_0110111011011100;
      90 : {coef1[11:0], coef0[18:0]} =   31'b110_100101111___001_0111000001101011;
      91 : {coef1[11:0], coef0[18:0]} =   31'b110_100101011___001_0111000111110101;
      92 : {coef1[11:0], coef0[18:0]} =   31'b110_100100111___001_0111001101111001;
      93 : {coef1[11:0], coef0[18:0]} =   31'b110_100100011___001_0111010011111000;
      94 : {coef1[11:0], coef0[18:0]} =   31'b110_100011111___001_0111011001110000;
      95 : {coef1[11:0], coef0[18:0]} =   31'b110_100011011___001_0111011111100001;
      96 : {coef1[11:0], coef0[18:0]} =   31'b110_100010111___001_0111100101001100;
      97 : {coef1[11:0], coef0[18:0]} =   31'b110_100010011___001_0111101010101111;
      98 : {coef1[11:0], coef0[18:0]} =   31'b110_100010000___001_0111110000001011;
      99 : {coef1[11:0], coef0[18:0]} =   31'b110_100001100___001_0111110101100000;
     100 : {coef1[11:0], coef0[18:0]} =   31'b110_100001001___001_0111111010101100;
     101 : {coef1[11:0], coef0[18:0]} =   31'b110_100000110___001_0111111111110001;
     102 : {coef1[11:0], coef0[18:0]} =   31'b110_100000011___001_1000000100101100;
     103 : {coef1[11:0], coef0[18:0]} =   31'b110_100000000___001_1000001001011111;
     104 : {coef1[11:0], coef0[18:0]} =   31'b110_011111101___001_1000001110001001;
     105 : {coef1[11:0], coef0[18:0]} =   31'b110_011111010___001_1000010010101010;
     106 : {coef1[11:0], coef0[18:0]} =   31'b110_011111000___001_1000010111000001;
     107 : {coef1[11:0], coef0[18:0]} =   31'b110_011110101___001_1000011011001110;
     108 : {coef1[11:0], coef0[18:0]} =   31'b110_011110011___001_1000011111010001;
     109 : {coef1[11:0], coef0[18:0]} =   31'b110_011110000___001_1000100011001010;
     110 : {coef1[11:0], coef0[18:0]} =   31'b110_011101110___001_1000100110111000;
     111 : {coef1[11:0], coef0[18:0]} =   31'b110_011101100___001_1000101010011011;
     112 : {coef1[11:0], coef0[18:0]} =   31'b110_011101010___001_1000101101110011;
     113 : {coef1[11:0], coef0[18:0]} =   31'b110_011101000___001_1000110000111111;
     114 : {coef1[11:0], coef0[18:0]} =   31'b110_011100111___001_1000110011111111;
     115 : {coef1[11:0], coef0[18:0]} =   31'b110_011100101___001_1000110110110100;
     116 : {coef1[11:0], coef0[18:0]} =   31'b110_011100100___001_1000111001011100;
     117 : {coef1[11:0], coef0[18:0]} =   31'b110_011100010___001_1000111011110111;
     118 : {coef1[11:0], coef0[18:0]} =   31'b110_011100001___001_1000111110000110;
     119 : {coef1[11:0], coef0[18:0]} =   31'b110_011100000___001_1001000000000111;
     120 : {coef1[11:0], coef0[18:0]} =   31'b110_011011111___001_1001000001111011;
     121 : {coef1[11:0], coef0[18:0]} =   31'b110_011011110___001_1001000011100010;
     122 : {coef1[11:0], coef0[18:0]} =   31'b110_011011110___001_1001000100111011;
     123 : {coef1[11:0], coef0[18:0]} =   31'b110_011011101___001_1001000110000101;
     124 : {coef1[11:0], coef0[18:0]} =   31'b110_011011101___001_1001000111000001;
     125 : {coef1[11:0], coef0[18:0]} =   31'b110_011011100___001_1001000111101111;
     126 : {coef1[11:0], coef0[18:0]} =   31'b110_011011100___001_1001001000001110;
     127 : {coef1[11:0], coef0[18:0]} =   31'b110_011011100___001_1001001000011101;
  endcase
end

endmodule // sin_cos_coef
